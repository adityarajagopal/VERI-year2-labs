library verilog;
use verilog.vl_types.all;
entity top is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end top;
